library verilog;
use verilog.vl_types.all;
entity Sea_Battle_vlg_vec_tst is
end Sea_Battle_vlg_vec_tst;
